LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Timer8254_tb IS
END Timer8254_tb;

ARCHITECTURE Behavioral OF Timer8254_tb IS

	COMPONENT Timer8254
		GENERIC (size : INTEGER);
		PORT (
			barcode_in : IN std_logic;
			clk : IN std_logic;
			en : IN std_logic;
			DACK : IN std_logic;
			rst : IN std_logic;
			captured_width : OUT std_logic_vector(size - 1 DOWNTO 0);
			DREQ : OUT std_logic);
	END COMPONENT;

	SIGNAL size : INTEGER := 16;
	SIGNAL barcode_in, DACK, clk, en, rst, DREQ : std_logic;
	SIGNAL captured_width : std_logic_vector(size - 1 DOWNTO 0);

BEGIN
	dut : Timer8254
	GENERIC MAP(size => size)
	PORT MAP(barcode_in => barcode_in, clk => clk, en => en, DACK => DACK, rst => rst, captured_width => captured_width, DREQ => DREQ);

	-- Clock process definitions
	clock_process : PROCESS
	BEGIN
		clk <= '0';
		WAIT FOR 25 ns;
		clk <= '1';
		WAIT FOR 25 ns;
	END PROCESS;

	handshake : PROCESS BEGIN
		IF (DREQ = '1') THEN
			DACK <= '1';
		ELSE
			DACK <= '0';
		END IF;
		WAIT FOR 100 ns;
	END PROCESS;
	-- Stimulus process
	stim_proc : PROCESS
	BEGIN
		barcode_in <= '1';
		rst <= '1';
		en <= '1';
		WAIT FOR 100 ns;
		rst <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		en <= '0';
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		en <= '1';
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		rst <= '1';
		barcode_in <= '0';
		WAIT FOR 200ns;
		rst <= '0';
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '0';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';
		WAIT FOR 200ns;
		barcode_in <= '1';

		WAIT;
	END PROCESS;
END Behavioral;